//this file is created for testing git functionality
//to be removed