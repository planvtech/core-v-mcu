module a2_bootrom
 #(
 parameter ADDR_WIDTH=32,
 parameter DATA_WIDTH=32
 )
 (
 input logic 		  CLK,
 input logic 		  CEN,
 input logic [ADDR_WIDTH-1:0]  A,
 output logic [DATA_WIDTH-1:0] Q
 );
 logic [31:0] 		  value;
 assign Q = value;
 always @(posedge CLK) begin
  case (A)
  0: value <= 32'h0B00006F;
  1: value <= 32'h0AC0006F;
  2: value <= 32'h0A80006F;
  3: value <= 32'h0A40006F;
  4: value <= 32'h0A00006F;
  5: value <= 32'h09C0006F;
  6: value <= 32'h0980006F;
  7: value <= 32'h0940006F;
  8: value <= 32'h0900006F;
  9: value <= 32'h08C0006F;
  10: value <= 32'h0880006F;
  11: value <= 32'h0840006F;
  12: value <= 32'h0800006F;
  13: value <= 32'h07C0006F;
  14: value <= 32'h0780006F;
  15: value <= 32'h0740006F;
  16: value <= 32'h0700006F;
  17: value <= 32'h06C0006F;
  18: value <= 32'h0680006F;
  19: value <= 32'h0640006F;
  20: value <= 32'h0600006F;
  21: value <= 32'h05C0006F;
  22: value <= 32'h0580006F;
  23: value <= 32'h0540006F;
  24: value <= 32'h0500006F;
  25: value <= 32'h04C0006F;
  26: value <= 32'h0480006F;
  27: value <= 32'h0440006F;
  28: value <= 32'h0400006F;
  29: value <= 32'h03C0006F;
  30: value <= 32'h0380006F;
  31: value <= 32'h0340006F;
  32: value <= 32'h0207C297;
  33: value <= 32'hF8028293;
  34: value <= 32'h0207E317;
  35: value <= 32'hF0030313;
  36: value <= 32'h0002A023;
  37: value <= 32'h00428293;
  38: value <= 32'hFE62ECE3;
  39: value <= 32'h0207E117;
  40: value <= 32'h2EC10113;
  41: value <= 32'h2270006F;
  42: value <= 32'h00060113;
  43: value <= 32'h00058067;
  44: value <= 32'h30200073;
  45: value <= 32'hC84A1101;
  46: value <= 32'h1C07E937;
  47: value <= 32'h4983C64E;
  48: value <= 32'hCC22F689;
  49: value <= 32'hCA26CE06;
  50: value <= 32'h842A4785;
  51: value <= 32'h06F98563;
  52: value <= 32'h00144783;
  53: value <= 32'h00044703;
  54: value <= 32'h8FD907A2;
  55: value <= 32'h07136729;
  56: value <= 32'h93635077;
  57: value <= 32'h478304E7;
  58: value <= 32'h07130064;
  59: value <= 32'h92630240;
  60: value <= 32'h470308E7;
  61: value <= 32'h47830034;
  62: value <= 32'h45030024;
  63: value <= 32'h07220054;
  64: value <= 32'h47838F5D;
  65: value <= 32'h46030044;
  66: value <= 32'h05620074;
  67: value <= 32'h8FD907C2;
  68: value <= 32'h00840593;
  69: value <= 32'h00EF8D5D;
  70: value <= 32'h47037550;
  71: value <= 32'h4785F689;
  72: value <= 32'h03100513;
  73: value <= 32'h02F70F63;
  74: value <= 32'h446240F2;
  75: value <= 32'h494244D2;
  76: value <= 32'h610549B2;
  77: value <= 32'h84AE8082;
  78: value <= 32'h05C215F9;
  79: value <= 32'h2D2D81C1;
  80: value <= 32'hC70394A2;
  81: value <= 32'hC783FFE4;
  82: value <= 32'h0722FFF4;
  83: value <= 32'h07C28FD9;
  84: value <= 32'h8FE383C1;
  85: value <= 32'h4783F6A7;
  86: value <= 32'h97E3F689;
  87: value <= 32'h0513FD37;
  88: value <= 32'h44620300;
  89: value <= 32'h44D240F2;
  90: value <= 32'h49B24942;
  91: value <= 32'h006F6105;
  92: value <= 32'h07137820;
  93: value <= 32'h92E30260;
  94: value <= 32'h1537FAE7;
  95: value <= 32'h05131A00;
  96: value <= 32'h259D1B05;
  97: value <= 32'h00344703;
  98: value <= 32'h00244783;
  99: value <= 32'h00544503;
  100: value <= 32'h8F5D0722;
  101: value <= 32'h00444783;
  102: value <= 32'h07C20562;
  103: value <= 32'h8D5D8FD9;
  104: value <= 32'h15372D55;
  105: value <= 32'h05131A00;
  106: value <= 32'h2D3D1E45;
  107: value <= 32'h00344783;
  108: value <= 32'h00244703;
  109: value <= 32'h8FD907A2;
  110: value <= 32'h00444703;
  111: value <= 32'h8F5D0742;
  112: value <= 32'h00544783;
  113: value <= 32'h8FD907E2;
  114: value <= 32'hA0019782;
  115: value <= 32'hC6061141;
  116: value <= 32'hC226C422;
  117: value <= 32'h00EFC04A;
  118: value <= 32'hC15170E0;
  119: value <= 32'hE7B74405;
  120: value <= 32'h80A31C07;
  121: value <= 32'hE7B7F887;
  122: value <= 32'h80231C07;
  123: value <= 32'h25EDF887;
  124: value <= 32'h1E6347E5;
  125: value <= 32'hE7B700F5;
  126: value <= 32'h84231C07;
  127: value <= 32'h4422F607;
  128: value <= 32'h449240B2;
  129: value <= 32'h05134902;
  130: value <= 32'h01410210;
  131: value <= 32'h25E9A5D5;
  132: value <= 32'h02000793;
  133: value <= 32'h00F51763;
  134: value <= 32'h1C07E7B7;
  135: value <= 32'hF6878423;
  136: value <= 32'h2D5DBFF9;
  137: value <= 32'h02300793;
  138: value <= 32'h02F51B63;
  139: value <= 32'h1C07E4B7;
  140: value <= 32'h89134401;
  141: value <= 32'hA8099284;
  142: value <= 32'h07B32551;
  143: value <= 32'h04050089;
  144: value <= 32'h80230442;
  145: value <= 32'h804100A7;
  146: value <= 32'hF57D2549;
  147: value <= 32'h442285A2;
  148: value <= 32'h490240B2;
  149: value <= 32'h92848513;
  150: value <= 32'h01414492;
  151: value <= 32'h40B2BDA1;
  152: value <= 32'h44924422;
  153: value <= 32'h01414902;
  154: value <= 32'h11018082;
  155: value <= 32'hCE06CA26;
  156: value <= 32'hC84ACC22;
  157: value <= 32'hC5194481;
  158: value <= 32'h84AE842A;
  159: value <= 32'h00B50933;
  160: value <= 32'h01241963;
  161: value <= 32'h446240F2;
  162: value <= 32'h85264942;
  163: value <= 32'h610544D2;
  164: value <= 32'h47838082;
  165: value <= 32'h06130004;
  166: value <= 32'h458500F1;
  167: value <= 32'h07A34501;
  168: value <= 32'h040500F1;
  169: value <= 32'h4E5000EF;
  170: value <= 32'h1537BFE1;
  171: value <= 32'h45911A00;
  172: value <= 32'h1D050513;
  173: value <= 32'h1537BF5D;
  174: value <= 32'h45AD1A00;
  175: value <= 32'h1C050513;
  176: value <= 32'h4785B76D;
  177: value <= 32'h00F51363;
  178: value <= 32'hE519B7CD;
  179: value <= 32'h1A001537;
  180: value <= 32'h051345A1;
  181: value <= 32'hBF511CC5;
  182: value <= 32'h80824501;
  183: value <= 32'hD4227179;
  184: value <= 32'h1C07E437;
  185: value <= 32'hF7D44783;
  186: value <= 32'hD226D606;
  187: value <= 32'hCE4ED04A;
  188: value <= 32'h000107A3;
  189: value <= 32'h6A634719;
  190: value <= 32'h173704F7;
  191: value <= 32'h078A1A00;
  192: value <= 32'h1F870713;
  193: value <= 32'h439C97BA;
  194: value <= 32'h00F10613;
  195: value <= 32'h45014585;
  196: value <= 32'h00EF8782;
  197: value <= 32'h47854AD0;
  198: value <= 32'h02F51963;
  199: value <= 32'h00F14703;
  200: value <= 32'h05300793;
  201: value <= 32'h02F71363;
  202: value <= 32'h1C07E7B7;
  203: value <= 32'hF817C703;
  204: value <= 32'hF6A40EA3;
  205: value <= 32'h80A3E319;
  206: value <= 32'hE7B7F8A7;
  207: value <= 32'hC7031C07;
  208: value <= 32'hE701F697;
  209: value <= 32'h84A34705;
  210: value <= 32'h50B2F6E7;
  211: value <= 32'h54925422;
  212: value <= 32'h49F25902;
  213: value <= 32'h80826145;
  214: value <= 32'h467000EF;
  215: value <= 32'h16E34785;
  216: value <= 32'h4783FEF5;
  217: value <= 32'hE73700F1;
  218: value <= 32'h0E231C07;
  219: value <= 32'h0713F6F7;
  220: value <= 32'h92630300;
  221: value <= 32'h478902E7;
  222: value <= 32'h1C07E737;
  223: value <= 32'hF6F71A23;
  224: value <= 32'hF6F40EA3;
  225: value <= 32'h1C07E7B7;
  226: value <= 32'hF6079F23;
  227: value <= 32'h1C07E7B7;
  228: value <= 32'hF6079523;
  229: value <= 32'h8793BF5D;
  230: value <= 32'hF793FCF7;
  231: value <= 32'h47210FF7;
  232: value <= 32'hFAF765E3;
  233: value <= 32'h1A001737;
  234: value <= 32'h0713078A;
  235: value <= 32'h97BA2147;
  236: value <= 32'h8782439C;
  237: value <= 32'h1C07E7B7;
  238: value <= 32'h9A23470D;
  239: value <= 32'h4789F6E7;
  240: value <= 32'hE7B7B7C1;
  241: value <= 32'h47111C07;
  242: value <= 32'h00EFBFCD;
  243: value <= 32'h47853F50;
  244: value <= 32'hF6F51DE3;
  245: value <= 32'h1C07E4B7;
  246: value <= 32'hF7E4D583;
  247: value <= 32'h00F14603;
  248: value <= 32'h1C07E6B7;
  249: value <= 32'hB2868713;
  250: value <= 32'h00B707B3;
  251: value <= 32'h00C78023;
  252: value <= 32'h00158793;
  253: value <= 32'h83C107C2;
  254: value <= 32'h00F56563;
  255: value <= 32'hF6F49F23;
  256: value <= 32'h0589B7A9;
  257: value <= 32'h05C2973E;
  258: value <= 32'h002381C1;
  259: value <= 32'h85130007;
  260: value <= 32'h9F23B286;
  261: value <= 32'h2515F6B4;
  262: value <= 32'h1C07E7B7;
  263: value <= 32'hF747D783;
  264: value <= 32'h81410542;
  265: value <= 32'h40F507B3;
  266: value <= 32'hE73717FD;
  267: value <= 32'h19231C07;
  268: value <= 32'hE7B7F6F7;
  269: value <= 32'hD7031C07;
  270: value <= 32'h9F23F6A7;
  271: value <= 32'h953AF604;
  272: value <= 32'hF6A79523;
  273: value <= 32'h0EA3478D;
  274: value <= 32'hB701F6F4;
  275: value <= 32'h373000EF;
  276: value <= 32'h1CE34785;
  277: value <= 32'hE4B7EEF5;
  278: value <= 32'hD5831C07;
  279: value <= 32'h4683F7E4;
  280: value <= 32'hE53700F1;
  281: value <= 32'h07131C07;
  282: value <= 32'h07B3B285;
  283: value <= 32'h802300B7;
  284: value <= 32'hE6B700D7;
  285: value <= 32'hD6831C07;
  286: value <= 32'h8793F746;
  287: value <= 32'h07C20015;
  288: value <= 32'h9F2383C1;
  289: value <= 32'h0686F6F4;
  290: value <= 32'hECD7C1E3;
  291: value <= 32'h973E0589;
  292: value <= 32'h81C105C2;
  293: value <= 32'h00070023;
  294: value <= 32'hB2850513;
  295: value <= 32'hF6B49F23;
  296: value <= 32'hE7B72B69;
  297: value <= 32'hE6B71C07;
  298: value <= 32'h57131C07;
  299: value <= 32'hAC230185;
  300: value <= 32'h7793F6A7;
  301: value <= 32'h97BA0FF5;
  302: value <= 32'hF6A6D703;
  303: value <= 32'hF6049F23;
  304: value <= 32'h571397BA;
  305: value <= 32'h77130085;
  306: value <= 32'h81410FF7;
  307: value <= 32'h751397BA;
  308: value <= 32'h97AA0FF5;
  309: value <= 32'hF6F69523;
  310: value <= 32'h1C07E7B7;
  311: value <= 32'hF6079723;
  312: value <= 32'h1C07E7B7;
  313: value <= 32'hF6079823;
  314: value <= 32'h1C07E7B7;
  315: value <= 32'hF7C7C783;
  316: value <= 32'h8713468D;
  317: value <= 32'h7713FD07;
  318: value <= 32'hE4630FF7;
  319: value <= 32'h479100E6;
  320: value <= 32'h8793B799;
  321: value <= 32'hF793FC97;
  322: value <= 32'h47090FF7;
  323: value <= 32'hE2F76FE3;
  324: value <= 32'hBF154795;
  325: value <= 32'h2AB000EF;
  326: value <= 32'h18E34785;
  327: value <= 32'hE4B7E2F5;
  328: value <= 32'hD7831C07;
  329: value <= 32'hE537F7E4;
  330: value <= 32'h46031C07;
  331: value <= 32'h071300F1;
  332: value <= 32'h06B3B285;
  333: value <= 32'h078500F7;
  334: value <= 32'h802307C2;
  335: value <= 32'h83C100C6;
  336: value <= 32'h9B634689;
  337: value <= 32'h478D02D7;
  338: value <= 32'h00070123;
  339: value <= 32'h0513458D;
  340: value <= 32'h9F23B285;
  341: value <= 32'h21D5F6F4;
  342: value <= 32'h1C07E7B7;
  343: value <= 32'hF707D703;
  344: value <= 32'h00170693;
  345: value <= 32'hF6D79823;
  346: value <= 32'h1C07E7B7;
  347: value <= 32'hA2878793;
  348: value <= 32'h802397BA;
  349: value <= 32'h478100A7;
  350: value <= 32'h1C07E6B7;
  351: value <= 32'hF6F49F23;
  352: value <= 32'hF6E6D783;
  353: value <= 32'h1C07E737;
  354: value <= 32'hF7275703;
  355: value <= 32'h07C20785;
  356: value <= 32'h972383C1;
  357: value <= 32'h0706F6F6;
  358: value <= 32'hDAE7C9E3;
  359: value <= 32'h1C07E5B7;
  360: value <= 32'hF6A5D703;
  361: value <= 32'h1C07E7B7;
  362: value <= 32'h1C07E637;
  363: value <= 32'hF707D803;
  364: value <= 32'h47814501;
  365: value <= 32'hA2860613;
  366: value <= 32'h0107EA63;
  367: value <= 32'h9523C119;
  368: value <= 32'h9F23F6E5;
  369: value <= 32'h9723F604;
  370: value <= 32'hB799F606;
  371: value <= 32'h00F60533;
  372: value <= 32'h00054503;
  373: value <= 32'hF7930785;
  374: value <= 32'h972A0FF7;
  375: value <= 32'h83410742;
  376: value <= 32'hBFD94505;
  377: value <= 32'h1DB000EF;
  378: value <= 32'h10E34785;
  379: value <= 32'hE4B7D6F5;
  380: value <= 32'hD5831C07;
  381: value <= 32'h4603F7E4;
  382: value <= 32'hE6B700F1;
  383: value <= 32'h87131C07;
  384: value <= 32'h07B3B286;
  385: value <= 32'h802300B7;
  386: value <= 32'h879300C7;
  387: value <= 32'h07C20015;
  388: value <= 32'h75E383C1;
  389: value <= 32'h0589DEF5;
  390: value <= 32'h05C2973E;
  391: value <= 32'h002381C1;
  392: value <= 32'h85130007;
  393: value <= 32'hE937B286;
  394: value <= 32'h9F231C07;
  395: value <= 32'h2131F6B4;
  396: value <= 32'hF6A95783;
  397: value <= 32'h0FF57513;
  398: value <= 32'h1C07E9B7;
  399: value <= 32'hFFF7C793;
  400: value <= 32'h0FF7F793;
  401: value <= 32'hF6A98623;
  402: value <= 32'hF6F91523;
  403: value <= 32'h06A79C63;
  404: value <= 32'h1C07E937;
  405: value <= 32'hF7892503;
  406: value <= 32'hE7B7C515;
  407: value <= 32'hC7831C07;
  408: value <= 32'h4689F7C7;
  409: value <= 32'hFCF78713;
  410: value <= 32'h0FF77713;
  411: value <= 32'h02E6E563;
  412: value <= 32'h1C07E7B7;
  413: value <= 32'hF707D603;
  414: value <= 32'h1C07E5B7;
  415: value <= 32'hA2858593;
  416: value <= 32'h1EB000EF;
  417: value <= 32'hE7B7311D;
  418: value <= 32'h98231C07;
  419: value <= 32'h9F23F607;
  420: value <= 32'h4799F604;
  421: value <= 32'h8793BB4D;
  422: value <= 32'hF793FC97;
  423: value <= 32'hE3E30FF7;
  424: value <= 32'h1537FEF6;
  425: value <= 32'h05131A00;
  426: value <= 32'h2A3D1D85;
  427: value <= 32'hF7892503;
  428: value <= 32'h15372255;
  429: value <= 32'h05131A00;
  430: value <= 32'h223D1E45;
  431: value <= 32'hF7892783;
  432: value <= 32'hA0019782;
  433: value <= 32'h1A001537;
  434: value <= 32'h1E850513;
  435: value <= 32'h55032A31;
  436: value <= 32'h2A0DF6A9;
  437: value <= 32'hF6C9C503;
  438: value <= 32'h45012235;
  439: value <= 32'hB76536DD;
  440: value <= 32'h0DF000EF;
  441: value <= 32'h12E34785;
  442: value <= 32'hE7B7C6F5;
  443: value <= 32'h8E231C07;
  444: value <= 32'hE7B7F607;
  445: value <= 32'hAC231C07;
  446: value <= 32'hE7B7F607;
  447: value <= 32'h97231C07;
  448: value <= 32'hE7B7F607;
  449: value <= 32'h9A231C07;
  450: value <= 32'hE7B7F607;
  451: value <= 32'h95231C07;
  452: value <= 32'hE7B7F607;
  453: value <= 32'h86231C07;
  454: value <= 32'hE7B7F607;
  455: value <= 32'h9F231C07;
  456: value <= 32'hE7B7F607;
  457: value <= 32'h98231C07;
  458: value <= 32'h0EA3F607;
  459: value <= 32'hB931F604;
  460: value <= 32'h1C07E737;
  461: value <= 32'h07136585;
  462: value <= 32'h4601D287;
  463: value <= 32'h02158593;
  464: value <= 32'h10000513;
  465: value <= 32'h00861793;
  466: value <= 32'h83C107C2;
  467: value <= 32'h981346A1;
  468: value <= 32'h58130107;
  469: value <= 32'h07864108;
  470: value <= 32'h00085363;
  471: value <= 32'h16FD8FAD;
  472: value <= 32'hF69307C2;
  473: value <= 32'h83C10FF6;
  474: value <= 32'h1023F2FD;
  475: value <= 32'h060500F7;
  476: value <= 32'h19E30709;
  477: value <= 32'h8082FCA6;
  478: value <= 32'hE63767C1;
  479: value <= 32'h86AA1C07;
  480: value <= 32'h85134701;
  481: value <= 32'h0613FFF7;
  482: value <= 32'h4363D286;
  483: value <= 32'h808200B7;
  484: value <= 32'h00E68833;
  485: value <= 32'h00084803;
  486: value <= 32'h00855793;
  487: value <= 32'hC7B30705;
  488: value <= 32'h07860107;
  489: value <= 32'hD80397B2;
  490: value <= 32'h17930007;
  491: value <= 32'h07C20085;
  492: value <= 32'h453383C1;
  493: value <= 32'hBFD100F8;
  494: value <= 32'hC62A1101;
  495: value <= 32'h45850070;
  496: value <= 32'hCE064505;
  497: value <= 32'h7C4000EF;
  498: value <= 32'h610540F2;
  499: value <= 32'h11418082;
  500: value <= 32'hC6064535;
  501: value <= 32'h40B237D5;
  502: value <= 32'h01414529;
  503: value <= 32'h47A9BFF1;
  504: value <= 32'h00F51363;
  505: value <= 32'hBFC9B7ED;
  506: value <= 32'hC4221141;
  507: value <= 32'h842AC606;
  508: value <= 32'h00040503;
  509: value <= 32'h40B2E509;
  510: value <= 32'h01414422;
  511: value <= 32'h37C58082;
  512: value <= 32'hB7FD0405;
  513: value <= 32'h00455793;
  514: value <= 32'h8BBD1141;
  515: value <= 32'hC606C422;
  516: value <= 32'h0713842A;
  517: value <= 32'h85130390;
  518: value <= 32'h54630307;
  519: value <= 32'h851300A7;
  520: value <= 32'h3F750577;
  521: value <= 32'h0513883D;
  522: value <= 32'h07930304;
  523: value <= 32'hD4630390;
  524: value <= 32'h051300A7;
  525: value <= 32'h44220574;
  526: value <= 32'h014140B2;
  527: value <= 32'h1141B74D;
  528: value <= 32'h842AC422;
  529: value <= 32'hC6068121;
  530: value <= 32'h85223F75;
  531: value <= 32'h40B24422;
  532: value <= 32'hBF4D0141;
  533: value <= 32'hC4221141;
  534: value <= 32'h8141842A;
  535: value <= 32'h37C5C606;
  536: value <= 32'h44228522;
  537: value <= 32'h014140B2;
  538: value <= 32'h77B7BFD9;
  539: value <= 32'h43881A10;
  540: value <= 32'h07F57513;
  541: value <= 32'h77378082;
  542: value <= 32'h47831A10;
  543: value <= 32'h75130007;
  544: value <= 32'hF79307F5;
  545: value <= 32'h8FC9F807;
  546: value <= 32'h00F70023;
  547: value <= 32'h47858082;
  548: value <= 32'h00F51F63;
  549: value <= 32'h1A107737;
  550: value <= 32'h00474783;
  551: value <= 32'h0017E793;
  552: value <= 32'h00F70223;
  553: value <= 32'h1A1077B7;
  554: value <= 32'h890543C8;
  555: value <= 32'hF97D8082;
  556: value <= 32'h1A107737;
  557: value <= 32'h00474783;
  558: value <= 32'hB7DD9BF9;
  559: value <= 32'h1A1077B7;
  560: value <= 32'h0847A503;
  561: value <= 32'h0FF57513;
  562: value <= 32'h77B78082;
  563: value <= 32'hA5031A10;
  564: value <= 32'h75130907;
  565: value <= 32'h80820FF5;
  566: value <= 32'h1A1077B7;
  567: value <= 32'h751343A8;
  568: value <= 32'h80820FF5;
  569: value <= 32'h1A1077B7;
  570: value <= 32'h751343E8;
  571: value <= 32'h80820FF5;
  572: value <= 32'h1A1077B7;
  573: value <= 32'h8082C7A8;
  574: value <= 32'hC2261141;
  575: value <= 32'h85936485;
  576: value <= 32'hC4224084;
  577: value <= 32'h842A4641;
  578: value <= 32'h450195AA;
  579: value <= 32'h94A2C606;
  580: value <= 32'hA60323AD;
  581: value <= 32'h47BD40C4;
  582: value <= 32'h02C7C063;
  583: value <= 32'h6585C205;
  584: value <= 32'h41858593;
  585: value <= 32'h442295A2;
  586: value <= 32'h449240B2;
  587: value <= 32'h06420612;
  588: value <= 32'h45418241;
  589: value <= 32'hA3910141;
  590: value <= 32'hB7D54641;
  591: value <= 32'h442240B2;
  592: value <= 32'h01414492;
  593: value <= 32'h71398082;
  594: value <= 32'h6985D64E;
  595: value <= 32'hD84ADC22;
  596: value <= 32'h892ACE5E;
  597: value <= 32'h41898413;
  598: value <= 32'hD2566B89;
  599: value <= 32'hDE06C66E;
  600: value <= 32'hD452DA26;
  601: value <= 32'hCC62D05A;
  602: value <= 32'hC86ACA66;
  603: value <= 32'h3769944A;
  604: value <= 32'h99CA4A81;
  605: value <= 32'h0DB79BCA;
  606: value <= 32'hA7830100;
  607: value <= 32'hE36340C9;
  608: value <= 32'h153702FA;
  609: value <= 32'h05131A00;
  610: value <= 32'h3DB924C5;
  611: value <= 32'h4109A503;
  612: value <= 32'h153735D1;
  613: value <= 32'h05131A00;
  614: value <= 32'h35B91E45;
  615: value <= 32'h4109A783;
  616: value <= 32'hA0019782;
  617: value <= 32'h1A0017B7;
  618: value <= 32'h23878513;
  619: value <= 32'h85563D35;
  620: value <= 32'h17B73555;
  621: value <= 32'h85131A00;
  622: value <= 32'h353D2547;
  623: value <= 32'h0C374048;
  624: value <= 32'h4C81E400;
  625: value <= 32'h2A033D41;
  626: value <= 32'h2B030044;
  627: value <= 32'h2D030004;
  628: value <= 32'h9C520084;
  629: value <= 32'hE5634454;
  630: value <= 32'h0A8500DC;
  631: value <= 32'hBF710441;
  632: value <= 32'h920BA483;
  633: value <= 32'h009D7563;
  634: value <= 32'h003D0493;
  635: value <= 32'h961398F1;
  636: value <= 32'h82410104;
  637: value <= 32'h01BC7B63;
  638: value <= 32'h855A85D2;
  639: value <= 32'h9A2629BD;
  640: value <= 32'h0D339B26;
  641: value <= 32'h0C85409D;
  642: value <= 32'h85CAB7F1;
  643: value <= 32'h21B5855A;
  644: value <= 32'h85CA8626;
  645: value <= 32'h2D918552;
  646: value <= 32'h4789B7DD;
  647: value <= 32'h00A7EE63;
  648: value <= 32'h00D087B7;
  649: value <= 32'h0516953E;
  650: value <= 32'h0737411C;
  651: value <= 32'h8FD90008;
  652: value <= 32'h411CC11C;
  653: value <= 32'hC11C9BED;
  654: value <= 32'h882A8082;
  655: value <= 32'h46814701;
  656: value <= 32'h43254501;
  657: value <= 32'h17934895;
  658: value <= 32'h83C10107;
  659: value <= 32'h00B7F963;
  660: value <= 32'h00E807B3;
  661: value <= 32'h0007C783;
  662: value <= 32'h0DF7F613;
  663: value <= 32'h8082E211;
  664: value <= 32'hFD078613;
  665: value <= 32'h0FF67613;
  666: value <= 32'h02C37B63;
  667: value <= 32'hFBF78613;
  668: value <= 32'h0FF67613;
  669: value <= 32'h00C8EC63;
  670: value <= 32'hFC978793;
  671: value <= 32'h0FF7F693;
  672: value <= 32'h00451793;
  673: value <= 32'h00F68533;
  674: value <= 32'hBF750705;
  675: value <= 32'hF9F78613;
  676: value <= 32'h0FF67613;
  677: value <= 32'hFEC8E6E3;
  678: value <= 32'hFA978793;
  679: value <= 32'h86B2B7C5;
  680: value <= 32'h6799B7C5;
  681: value <= 32'h87931101;
  682: value <= 32'h16235487;
  683: value <= 32'h450100F1;
  684: value <= 32'h06C00793;
  685: value <= 32'h0723CE06;
  686: value <= 32'h231D00F1;
  687: value <= 32'h458D0070;
  688: value <= 32'h2B8D4501;
  689: value <= 32'h610540F2;
  690: value <= 32'h71398082;
  691: value <= 32'hDE064501;
  692: value <= 32'hDA26DC22;
  693: value <= 32'hD64ED84A;
  694: value <= 32'hCC02D452;
  695: value <= 32'h3F35CE02;
  696: value <= 32'h3F254505;
  697: value <= 32'h3F154509;
  698: value <= 32'h1A1047B7;
  699: value <= 32'h0D87A703;
  700: value <= 32'hCA3A4505;
  701: value <= 32'h0C47A703;
  702: value <= 32'hC63A8B05;
  703: value <= 32'h0C47A783;
  704: value <= 32'hC63E8B85;
  705: value <= 32'h33953369;
  706: value <= 32'h06200793;
  707: value <= 32'h00F50563;
  708: value <= 32'h06200513;
  709: value <= 32'h6471338D;
  710: value <= 32'h20040593;
  711: value <= 32'h21194501;
  712: value <= 32'h20040593;
  713: value <= 32'h2EFD4505;
  714: value <= 32'h15373FAD;
  715: value <= 32'h05131A00;
  716: value <= 32'h395D25C5;
  717: value <= 32'h1A001537;
  718: value <= 32'h26850513;
  719: value <= 32'h15373175;
  720: value <= 32'h05131A00;
  721: value <= 32'h314D26C5;
  722: value <= 32'h1A001537;
  723: value <= 32'h27850513;
  724: value <= 32'h47323961;
  725: value <= 32'h18634785;
  726: value <= 32'h15370CF7;
  727: value <= 32'h05131A00;
  728: value <= 32'h31592905;
  729: value <= 32'h1A001537;
  730: value <= 32'h29850513;
  731: value <= 32'h455239B5;
  732: value <= 32'h25B73951;
  733: value <= 32'h85930026;
  734: value <= 32'h45015A05;
  735: value <= 32'h458122BD;
  736: value <= 32'h24354501;
  737: value <= 32'h45014581;
  738: value <= 32'h45012471;
  739: value <= 32'h47852A59;
  740: value <= 32'h47B2C83E;
  741: value <= 32'h0793EFD1;
  742: value <= 32'h0C2302E0;
  743: value <= 32'h47B200F1;
  744: value <= 32'h00010CA3;
  745: value <= 32'h9E634705;
  746: value <= 32'h47420AE7;
  747: value <= 32'h0AF71B63;
  748: value <= 32'h1C07C537;
  749: value <= 32'h04136785;
  750: value <= 32'h64890005;
  751: value <= 32'h00940933;
  752: value <= 32'h00050513;
  753: value <= 32'h2023943E;
  754: value <= 32'h2E2392F9;
  755: value <= 32'h22239009;
  756: value <= 32'h22234004;
  757: value <= 32'h330D9209;
  758: value <= 32'h92092783;
  759: value <= 32'h40C42803;
  760: value <= 32'h1C07D737;
  761: value <= 32'hFFF78893;
  762: value <= 32'h40F006B3;
  763: value <= 32'h41C70713;
  764: value <= 32'h05374601;
  765: value <= 32'h84931C00;
  766: value <= 32'h10639284;
  767: value <= 32'h67890506;
  768: value <= 32'h660597AA;
  769: value <= 32'h92C7A023;
  770: value <= 32'h51960613;
  771: value <= 32'h15B7962A;
  772: value <= 32'hAE231A00;
  773: value <= 32'hA2239007;
  774: value <= 32'h06139207;
  775: value <= 32'h85934006;
  776: value <= 32'hF0EF9465;
  777: value <= 32'h1537C86F;
  778: value <= 32'h05131A00;
  779: value <= 32'hBF152945;
  780: value <= 32'hF7B547C2;
  781: value <= 32'h02100793;
  782: value <= 32'h431CB78D;
  783: value <= 32'h00F56963;
  784: value <= 32'h95BE434C;
  785: value <= 32'h00B56963;
  786: value <= 32'h07410605;
  787: value <= 32'h05B3B77D;
  788: value <= 32'hFBE30095;
  789: value <= 32'h434CFEB7;
  790: value <= 32'h97C697AE;
  791: value <= 32'h00D7F533;
  792: value <= 32'h34F9B7E5;
  793: value <= 32'h1A1047B7;
  794: value <= 32'hA683C602;
  795: value <= 32'h47050D87;
  796: value <= 32'h02700513;
  797: value <= 32'h00E68863;
  798: value <= 32'h0D87A783;
  799: value <= 32'hC7818B89;
  800: value <= 32'h02800513;
  801: value <= 32'h47B731B5;
  802: value <= 32'h47051A10;
  803: value <= 32'hDBF86459;
  804: value <= 32'h1A1044B7;
  805: value <= 32'h1C07E937;
  806: value <= 32'h1C07E9B7;
  807: value <= 32'hF8F40413;
  808: value <= 32'h58FC4A05;
  809: value <= 32'h01478863;
  810: value <= 32'h1C0087B7;
  811: value <= 32'h08078793;
  812: value <= 32'hA0019782;
  813: value <= 32'hF8094783;
  814: value <= 32'hF0EFE399;
  815: value <= 32'hC783E22F;
  816: value <= 32'hE399F699;
  817: value <= 32'hD08FF0EF;
  818: value <= 32'h078547B2;
  819: value <= 32'h47B2C63E;
  820: value <= 32'hFCF479E3;
  821: value <= 32'h1C07E7B7;
  822: value <= 32'hF817C783;
  823: value <= 32'h0828E789;
  824: value <= 32'hF0EF3621;
  825: value <= 32'hC602DD4F;
  826: value <= 32'h2737BF65;
  827: value <= 32'h47141A10;
  828: value <= 32'h95334791;
  829: value <= 32'h8EC900A7;
  830: value <= 32'h4714C714;
  831: value <= 32'hFFF54793;
  832: value <= 32'hC71C8FF5;
  833: value <= 32'h8D5D431C;
  834: value <= 32'h004C57B7;
  835: value <= 32'hB4078793;
  836: value <= 32'h02B7D7B3;
  837: value <= 32'hE737C308;
  838: value <= 32'h45011C07;
  839: value <= 32'hF8F70123;
  840: value <= 32'h27B78082;
  841: value <= 32'hC7031A10;
  842: value <= 32'hE6B71887;
  843: value <= 32'h87931C07;
  844: value <= 32'h9B3D1807;
  845: value <= 32'h00E78423;
  846: value <= 32'h0187C703;
  847: value <= 32'h8C239B3D;
  848: value <= 32'hC70300E7;
  849: value <= 32'h9B3D0287;
  850: value <= 32'h02E78423;
  851: value <= 32'hF826C683;
  852: value <= 32'h1C07E737;
  853: value <= 32'hF2D72423;
  854: value <= 32'hF2870713;
  855: value <= 32'h100006B7;
  856: value <= 32'h06B7C354;
  857: value <= 32'h86932007;
  858: value <= 32'hC71409F6;
  859: value <= 32'h704706B7;
  860: value <= 32'hC754068D;
  861: value <= 32'h900006B7;
  862: value <= 32'hCB140685;
  863: value <= 32'h4691C388;
  864: value <= 32'hC683C3D4;
  865: value <= 32'hE6930087;
  866: value <= 32'h84230106;
  867: value <= 32'hD39800D7;
  868: value <= 32'hD3D84751;
  869: value <= 32'h0287C703;
  870: value <= 32'h01076713;
  871: value <= 32'h02E78423;
  872: value <= 32'h1A102737;
  873: value <= 32'h18070793;
  874: value <= 32'hFFED43DC;
  875: value <= 32'h27B78082;
  876: value <= 32'h87930034;
  877: value <= 32'h953E0437;
  878: value <= 32'h4783051E;
  879: value <= 32'hE7370285;
  880: value <= 32'h47031C07;
  881: value <= 32'h9BBDF827;
  882: value <= 32'h02F50423;
  883: value <= 32'h02854783;
  884: value <= 32'h0407E793;
  885: value <= 32'h02F50423;
  886: value <= 32'h1C07E7B7;
  887: value <= 32'hF2E7A423;
  888: value <= 32'h10000737;
  889: value <= 32'h07378DD9;
  890: value <= 32'h87932007;
  891: value <= 32'h0713F287;
  892: value <= 32'hC7980667;
  893: value <= 32'h90000737;
  894: value <= 32'hD11C0705;
  895: value <= 32'hC7D8C3CC;
  896: value <= 32'hD15C47C1;
  897: value <= 32'h02854783;
  898: value <= 32'h0107E793;
  899: value <= 32'h02F50423;
  900: value <= 32'h80824501;
  901: value <= 32'h003427B7;
  902: value <= 32'h04378793;
  903: value <= 32'h051E953E;
  904: value <= 32'h02854783;
  905: value <= 32'h1C07E737;
  906: value <= 32'hF8274703;
  907: value <= 32'h04239BBD;
  908: value <= 32'h478302F5;
  909: value <= 32'hE7930285;
  910: value <= 32'h04230407;
  911: value <= 32'hE7B702F5;
  912: value <= 32'hA4231C07;
  913: value <= 32'h0737F2E7;
  914: value <= 32'h8DD91000;
  915: value <= 32'h20070737;
  916: value <= 32'hF2878793;
  917: value <= 32'h09970713;
  918: value <= 32'h0737C798;
  919: value <= 32'h07059000;
  920: value <= 32'hC3CCD11C;
  921: value <= 32'h47C1C7D8;
  922: value <= 32'h4783D15C;
  923: value <= 32'hE7930285;
  924: value <= 32'h04230107;
  925: value <= 32'h450102F5;
  926: value <= 32'h27B78082;
  927: value <= 32'hC7031A10;
  928: value <= 32'hE6B71887;
  929: value <= 32'h08371C07;
  930: value <= 32'h9B3D2007;
  931: value <= 32'h18E78423;
  932: value <= 32'h1987C703;
  933: value <= 32'h200F08B7;
  934: value <= 32'h18078793;
  935: value <= 32'h8C239B3D;
  936: value <= 32'hC70300E7;
  937: value <= 32'h9B3D0287;
  938: value <= 32'h02E78423;
  939: value <= 32'hF826C683;
  940: value <= 32'h1C07E737;
  941: value <= 32'hF2D72423;
  942: value <= 32'hF2870713;
  943: value <= 32'h100006B7;
  944: value <= 32'h0693C354;
  945: value <= 32'hC7140038;
  946: value <= 32'h00855693;
  947: value <= 32'h82C106C2;
  948: value <= 32'h0FF57513;
  949: value <= 32'h0116E6B3;
  950: value <= 32'h01056533;
  951: value <= 32'hCB08C754;
  952: value <= 32'hFFF60693;
  953: value <= 32'h70470537;
  954: value <= 32'hCB548EC9;
  955: value <= 32'h900006B7;
  956: value <= 32'hCF140685;
  957: value <= 32'hC3D0C38C;
  958: value <= 32'h0087C683;
  959: value <= 32'h0106E693;
  960: value <= 32'h00D78423;
  961: value <= 32'h4771D398;
  962: value <= 32'hC703D3D8;
  963: value <= 32'h67130287;
  964: value <= 32'h84230107;
  965: value <= 32'h273702E7;
  966: value <= 32'h07931A10;
  967: value <= 32'h43DC1807;
  968: value <= 32'h8082FFED;
  969: value <= 32'h1A102737;
  970: value <= 32'h47854714;
  971: value <= 32'h00A797B3;
  972: value <= 32'hC7148EDD;
  973: value <= 32'hC6934710;
  974: value <= 32'h8EF1FFF7;
  975: value <= 32'h4314C714;
  976: value <= 32'hC31C8FD5;
  977: value <= 32'h003427B7;
  978: value <= 32'h04178793;
  979: value <= 32'h57B7953E;
  980: value <= 32'h8793004C;
  981: value <= 32'hD7B3B407;
  982: value <= 32'h051E02B7;
  983: value <= 32'h83C107C2;
  984: value <= 32'h02F51323;
  985: value <= 32'hE793515C;
  986: value <= 32'hD15C0067;
  987: value <= 32'hE793515C;
  988: value <= 32'hD15C0107;
  989: value <= 32'hE793515C;
  990: value <= 32'hD15C1007;
  991: value <= 32'hE793515C;
  992: value <= 32'hD15C2007;
  993: value <= 32'h80824501;
  994: value <= 32'h003427B7;
  995: value <= 32'h04178793;
  996: value <= 32'h1793953E;
  997: value <= 32'h45010075;
  998: value <= 32'hEF114BD8;
  999: value <= 32'hCBCCCB90;
  1000: value <= 32'h0187C703;
  1001: value <= 32'h01076713;
  1002: value <= 32'h00E78C23;
  1003: value <= 32'hE7114BD8;
  1004: value <= 32'h81410542;
  1005: value <= 32'h05058082;
  1006: value <= 32'h0505B7C5;
  1007: value <= 32'h27B7BFC5;
  1008: value <= 32'h87930034;
  1009: value <= 32'h953E0417;
  1010: value <= 32'h591C051E;
  1011: value <= 32'hC7998B85;
  1012: value <= 32'h03454783;
  1013: value <= 32'h00234505;
  1014: value <= 32'h808200F6;
  1015: value <= 32'h80824501;
  1016: value <= 32'h1A102737;
  1017: value <= 32'h07934714;
  1018: value <= 32'h97B32000;
  1019: value <= 32'h8EDD00A7;
  1020: value <= 32'h4710C714;
  1021: value <= 32'hFFF7C693;
  1022: value <= 32'hC7148EF1;
  1023: value <= 32'h8FD54314;
  1024: value <= 32'h27B7C31C;
  1025: value <= 32'h87930034;
  1026: value <= 32'h953E04A7;
  1027: value <= 32'h5783051E;
  1028: value <= 32'hE79301C5;
  1029: value <= 32'h1E231007;
  1030: value <= 32'hE7B700F5;
  1031: value <= 32'hA7831C07;
  1032: value <= 32'hC11CF847;
  1033: value <= 32'h01C55783;
  1034: value <= 32'h2007E793;
  1035: value <= 32'h00F51E23;
  1036: value <= 32'h80824501;
  1037: value <= 32'h003427B7;
  1038: value <= 32'h04A78793;
  1039: value <= 32'h1793953E;
  1040: value <= 32'h45010075;
  1041: value <= 32'hEF114B98;
  1042: value <= 32'hCB8CC7D0;
  1043: value <= 32'h0147C703;
  1044: value <= 32'h01076713;
  1045: value <= 32'h00E78A23;
  1046: value <= 32'hE7114B98;
  1047: value <= 32'h81410542;
  1048: value <= 32'h05058082;
  1049: value <= 32'h0505B7C5;
  1050: value <= 32'h47B3BFC5;
  1051: value <= 32'h8B8D00B5;
  1052: value <= 32'h00C508B3;
  1053: value <= 32'h478DE7B1;
  1054: value <= 32'h04C7F463;
  1055: value <= 32'h00357793;
  1056: value <= 32'hEBB9872A;
  1057: value <= 32'hFFC8F613;
  1058: value <= 32'h40E606B3;
  1059: value <= 32'h02000793;
  1060: value <= 32'h06D7C863;
  1061: value <= 32'h87BA86AE;
  1062: value <= 32'h02C77163;
  1063: value <= 32'h0006A803;
  1064: value <= 32'h06910791;
  1065: value <= 32'hFF07AE23;
  1066: value <= 32'hFEC7EAE3;
  1067: value <= 32'hFFF60793;
  1068: value <= 32'h9BF18F99;
  1069: value <= 32'h973E0791;
  1070: value <= 32'h666395BE;
  1071: value <= 32'h80820117;
  1072: value <= 32'h7E63872A;
  1073: value <= 32'hC7830315;
  1074: value <= 32'h07050005;
  1075: value <= 32'h0FA30585;
  1076: value <= 32'h9AE3FEF7;
  1077: value <= 32'h8082FEE8;
  1078: value <= 32'h0005C683;
  1079: value <= 32'h77930705;
  1080: value <= 32'h0FA30037;
  1081: value <= 32'h0585FED7;
  1082: value <= 32'hC683DFD1;
  1083: value <= 32'h07050005;
  1084: value <= 32'h00377793;
  1085: value <= 32'hFED70FA3;
  1086: value <= 32'hFFF90585;
  1087: value <= 32'h8082B761;
  1088: value <= 32'hC6221141;
  1089: value <= 32'h02000413;
  1090: value <= 32'h0005A383;
  1091: value <= 32'h0045A283;
  1092: value <= 32'h0085AF83;
  1093: value <= 32'h00C5AF03;
  1094: value <= 32'h0105AE83;
  1095: value <= 32'h0145AE03;
  1096: value <= 32'h0185A303;
  1097: value <= 32'h01C5A803;
  1098: value <= 32'h07135194;
  1099: value <= 32'h07B30247;
  1100: value <= 32'h2E2340E6;
  1101: value <= 32'h2023FC77;
  1102: value <= 32'h2223FE57;
  1103: value <= 32'h2423FFF7;
  1104: value <= 32'h2623FFE7;
  1105: value <= 32'h2823FFD7;
  1106: value <= 32'h2A23FFC7;
  1107: value <= 32'h2C23FE67;
  1108: value <= 32'h2E23FF07;
  1109: value <= 32'h8593FED7;
  1110: value <= 32'h47E30245;
  1111: value <= 32'h86AEFAF4;
  1112: value <= 32'h716387BA;
  1113: value <= 32'hA80302C7;
  1114: value <= 32'h07910006;
  1115: value <= 32'hAE230691;
  1116: value <= 32'hEAE3FF07;
  1117: value <= 32'h0793FEC7;
  1118: value <= 32'h8F99FFF6;
  1119: value <= 32'h07919BF1;
  1120: value <= 32'h95BE973E;
  1121: value <= 32'h01176563;
  1122: value <= 32'h01414432;
  1123: value <= 32'hC7838082;
  1124: value <= 32'h07050005;
  1125: value <= 32'h0FA30585;
  1126: value <= 32'h87E3FEF7;
  1127: value <= 32'hC783FEE8;
  1128: value <= 32'h07050005;
  1129: value <= 32'h0FA30585;
  1130: value <= 32'h92E3FEF7;
  1131: value <= 32'hBFE9FEE8;
  1132: value <= 32'h4332490A;
  1133: value <= 32'h204C4220;
  1134: value <= 32'h20504D4A;
  1135: value <= 32'h00000000;
  1136: value <= 32'h42203241;
  1137: value <= 32'h4D544F4F;
  1138: value <= 32'h000A0D45;
  1139: value <= 32'h20544F4E;
  1140: value <= 32'h0A0D4B4F;
  1141: value <= 32'h00000000;
  1142: value <= 32'h5241550A;
  1143: value <= 32'h4C422054;
  1144: value <= 32'h504D4A20;
  1145: value <= 32'h00000020;
  1146: value <= 32'h4B48430A;
  1147: value <= 32'h204D5553;
  1148: value <= 32'h20525245;
  1149: value <= 32'h00000000;
  1150: value <= 32'h1A000312;
  1151: value <= 32'h1A000358;
  1152: value <= 32'h1A0003CA;
  1153: value <= 32'h1A00044C;
  1154: value <= 32'h1A000514;
  1155: value <= 32'h1A0005E4;
  1156: value <= 32'h1A0006E0;
  1157: value <= 32'h1A000376;
  1158: value <= 32'h1A0003B4;
  1159: value <= 32'h1A0003C2;
  1160: value <= 32'h1A00034A;
  1161: value <= 32'h1A0003BE;
  1162: value <= 32'h1A00034A;
  1163: value <= 32'h1A0003C2;
  1164: value <= 32'h1A0003B4;
  1165: value <= 32'h1A000376;
  1166: value <= 32'h616F4C0A;
  1167: value <= 32'h676E6964;
  1168: value <= 32'h63655320;
  1169: value <= 32'h6E6F6974;
  1170: value <= 32'h00000020;
  1171: value <= 32'h6D754A0A;
  1172: value <= 32'h676E6970;
  1173: value <= 32'h206F7420;
  1174: value <= 32'h00000000;
  1175: value <= 32'h2072614D;
  1176: value <= 32'h32203120;
  1177: value <= 32'h00333230;
  1178: value <= 32'h00002020;
  1179: value <= 32'h323A3931;
  1180: value <= 32'h31303A32;
  1181: value <= 32'h00000000;
  1182: value <= 32'h2032410A;
  1183: value <= 32'h746F6F42;
  1184: value <= 32'h64616F6C;
  1185: value <= 32'h42207265;
  1186: value <= 32'h73746F6F;
  1187: value <= 32'h003D6C65;
  1188: value <= 32'h00002031;
  1189: value <= 32'h00002030;
  1190: value <= 32'h003D7272;
  default: value <= 0;
   endcase
  end
endmodule    
